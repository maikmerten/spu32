// !!! IN MOST SITUATIONS YOU DO NOT NEED TO EDIT THIS FILE. !!!
//
// This file is a template for your local build config. The file config-local.vh
// is initially created from this template. Modify config-local.vh instead.
// Invoke 'make config-local.vh" and edit config-local.vh if you want to edit
// the system configuration.


// === Extension board configuration ===
// Uncomment the following define if you have the HX8K Breakout Board Extension.
// Information about that extension board:
//    https://github.com/maikmerten/hx8k-breakout-extension
// With the extension board present, RAM capacity is 512 KB.
// Without the extension board, RAM capacity is 8 KB.

//`define EXTENSION_PRESENT


// === Cache configuration ===
// Uncomment the following define if you want to include a CPU cache. This improves
// CPU perfomance by about 25%, but increases FPGA utilization a bit.

//`define ENABLE_CACHE
